  --Example instantiation for system 'mon_sopc'
  mon_sopc_inst : mon_sopc
    port map(
      ledBabord_from_the_avalon_Gestion_0 => ledBabord_from_the_avalon_Gestion_0,
      ledSTBY_from_the_avalon_Gestion_0 => ledSTBY_from_the_avalon_Gestion_0,
      ledTribord_from_the_avalon_Gestion_0 => ledTribord_from_the_avalon_Gestion_0,
      out_bip_from_the_avalon_Gestion_0 => out_bip_from_the_avalon_Gestion_0,
      BP_Babord_to_the_avalon_Gestion_0 => BP_Babord_to_the_avalon_Gestion_0,
      BP_STBY_to_the_avalon_Gestion_0 => BP_STBY_to_the_avalon_Gestion_0,
      BP_Tribord_to_the_avalon_Gestion_0 => BP_Tribord_to_the_avalon_Gestion_0,
      clk_0 => clk_0,
      reset_n => reset_n
    );


